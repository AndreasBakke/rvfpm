/*  rvfpm - 2024
  Andreas S. Bakke

  Description:
  RISC-V Floating Point Unit Model.
  Package for types
*/
`include "defines.svh"
package pa_rvfpm;

endpackage : pa_rvfpm

